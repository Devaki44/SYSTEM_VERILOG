//CODE
class packet #(int unsigned N = 31);
  rand bit[31:0] data;
  rand bit[31:0] k;

constraint power_of_two {k inside {[0:N]};        
                         data == (1 << k);}
endclass

module test;
  packet#(31) pkt;
  initial begin
    pkt = new();
    
    repeat(32)begin
      pkt.randomize();
      $display(" data = %b ",pkt.data);
    end
  end
endmodule


//OUTPUT
 data = 00000000000000000000010000000000 
 data = 00010000000000000000000000000000 
 data = 00000000000000000001000000000000 
 data = 00000010000000000000000000000000 
 data = 00000010000000000000000000000000 
 data = 10000000000000000000000000000000 
 data = 00000000000000100000000000000000 
 data = 10000000000000000000000000000000 
 data = 00000000001000000000000000000000 
 data = 00000000000000000000000000010000 
 data = 00000000000000000000000010000000 
 data = 00000000001000000000000000000000 
 data = 00000000000001000000000000000000 
 data = 00000000000000000000000000100000 
 data = 10000000000000000000000000000000 
 data = 00000000001000000000000000000000 
 data = 00000000000010000000000000000000 
 data = 00000000001000000000000000000000 
 data = 00000000000000000000000000010000 
 data = 00000000100000000000000000000000 
 data = 00000000000000000001000000000000 
 data = 00000000000000000000100000000000 
 data = 00000000000000000000000000000100 
 data = 00010000000000000000000000000000 
 data = 00000000000000000000000100000000 
 data = 00000000000000001000000000000000 
 data = 00000000010000000000000000000000 
 data = 00000000000000000000010000000000 
 data = 00000000000000000001000000000000 
 data = 00000000000000000000000100000000 
 data = 00000000000000000000000000001000 
 data = 00000100000000000000000000000000 
           V C S   S i m u l a t i o n   R e p o r t 
