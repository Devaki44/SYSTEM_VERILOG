
module Unpacked_array;
  byte a[7:0];
  
  initial begin
    
    foreach(a[i])begin
      
      a[i] = $urandom_range(0,64);
      
      $display("data of a[%0d] = %b",i,a[i]);
    end
  end
endmodule

# KERNEL: data of a[7] = 00101010
# KERNEL: data of a[6] = 00110100
# KERNEL: data of a[5] = 00101101
# KERNEL: data of a[4] = 00100100
# KERNEL: data of a[3] = 00010101
# KERNEL: data of a[2] = 00001011
# KERNEL: data of a[1] = 00001010
# KERNEL: data of a[0] = 01000000
# KERNEL: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.




module Unpacked_array;
  int a[31:0];
  
  initial begin
    
    foreach(a[i])begin
      
      a[i] = $urandom_range(0,4096);
      
      $display("data of a[%0d] = %b",i,a[i]);
    end
  end
endmodule

# KERNEL: data of a[31] = 00000000000000000000110101110101
# KERNEL: data of a[30] = 00000000000000000000011100011111
# KERNEL: data of a[29] = 00000000000000000000101110000010
# KERNEL: data of a[28] = 00000000000000000000100110001110
# KERNEL: data of a[27] = 00000000000000000000000011000001
# KERNEL: data of a[26] = 00000000000000000000000011100011
# KERNEL: data of a[25] = 00000000000000000000101101110110
# KERNEL: data of a[24] = 00000000000000000000111100110111
# KERNEL: data of a[23] = 00000000000000000000010100100010
# KERNEL: data of a[22] = 00000000000000000000011110110010
# KERNEL: data of a[21] = 00000000000000000000101011001010
# KERNEL: data of a[20] = 00000000000000000000101111010100
# KERNEL: data of a[19] = 00000000000000000000110011010010
# KERNEL: data of a[18] = 00000000000000000000111110101000
# KERNEL: data of a[17] = 00000000000000000000101000011101
# KERNEL: data of a[16] = 00000000000000000000001010000001
# KERNEL: data of a[15] = 00000000000000000000100100011111
# KERNEL: data of a[14] = 00000000000000000000001111010000
# KERNEL: data of a[13] = 00000000000000000000010101100001
# KERNEL: data of a[12] = 00000000000000000000100001100100
# KERNEL: data of a[11] = 00000000000000000000001111001101
# KERNEL: data of a[10] = 00000000000000000000101000101111
# KERNEL: data of a[9] = 00000000000000000000001001100001
# KERNEL: data of a[8] = 00000000000000000000001110100101
# KERNEL: data of a[7] = 00000000000000000000010001110100
# KERNEL: data of a[6] = 00000000000000000000011101010010
# KERNEL: data of a[5] = 00000000000000000000000101010100
# KERNEL: data of a[4] = 00000000000000000000000101110010
# KERNEL: data of a[3] = 00000000000000000000111110000011
# KERNEL: data of a[2] = 00000000000000000000110010111111
# KERNEL: data of a[1] = 00000000000000000000111000110110
# KERNEL: data of a[0] = 00000000000000000000100001101010
# KERNEL: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.




module Unpacked_array;
  shortint a[15:0];
  
  initial begin
    
    foreach(a[i])begin
      
      a[i] = $urandom_range(0,4096);
      
      $display("data of a[%0d] = %b",i,a[i]);
    end
  end
endmodule

# KERNEL: data of a[15] = 0000110101110101
# KERNEL: data of a[14] = 0000011100011111
# KERNEL: data of a[13] = 0000101110000010
# KERNEL: data of a[12] = 0000100110001110
# KERNEL: data of a[11] = 0000000011000001
# KERNEL: data of a[10] = 0000000011100011
# KERNEL: data of a[9] = 0000101101110110
# KERNEL: data of a[8] = 0000111100110111
# KERNEL: data of a[7] = 0000010100100010
# KERNEL: data of a[6] = 0000011110110010
# KERNEL: data of a[5] = 0000101011001010
# KERNEL: data of a[4] = 0000101111010100
# KERNEL: data of a[3] = 0000110011010010
# KERNEL: data of a[2] = 0000111110101000
# KERNEL: data of a[1] = 0000101000011101
# KERNEL: data of a[0] = 0000001010000001
# KERNEL: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.




module Unpacked_array;
  longint a[63:0];
  
  initial begin
    
    foreach(a[i])begin
      
      a[i] = $urandom_range(0,409600);
      
      $display("data of a[%0d] = %b",i,a[i]);
    end
  end
endmodule
# KERNEL: data of a[63] = 0000000000000000000000000000000000000000000001100000010011000010
# KERNEL: data of a[62] = 0000000000000000000000000000000000000000000001000000000011101011
# KERNEL: data of a[61] = 0000000000000000000000000000000000000000000001001010001111111100
# KERNEL: data of a[60] = 0000000000000000000000000000000000000000000000100000000010010010
# KERNEL: data of a[59] = 0000000000000000000000000000000000000000000001011100001100001010
# KERNEL: data of a[58] = 0000000000000000000000000000000000000000000000111010100011110101
# KERNEL: data of a[57] = 0000000000000000000000000000000000000000000000000001111000100100
# KERNEL: data of a[56] = 0000000000000000000000000000000000000000000000101011100001101011
# KERNEL: data of a[55] = 0000000000000000000000000000000000000000000001001100101100110000
# KERNEL: data of a[54] = 0000000000000000000000000000000000000000000001011010011100110101
# KERNEL: data of a[53] = 0000000000000000000000000000000000000000000000101011100110010111
# KERNEL: data of a[52] = 0000000000000000000000000000000000000000000001011001001101100000
# KERNEL: data of a[51] = 0000000000000000000000000000000000000000000001010001101001011000
# KERNEL: data of a[50] = 0000000000000000000000000000000000000000000000011110111101000111
# KERNEL: data of a[49] = 0000000000000000000000000000000000000000000000001110001010000101
# KERNEL: data of a[48] = 0000000000000000000000000000000000000000000000011110100010101110
# KERNEL: data of a[47] = 0000000000000000000000000000000000000000000000010101000001110100
# KERNEL: data of a[46] = 0000000000000000000000000000000000000000000001010001100100001111
# KERNEL: data of a[45] = 0000000000000000000000000000000000000000000001001100011111101000
# KERNEL: data of a[44] = 0000000000000000000000000000000000000000000000111111100111100011
# KERNEL: data of a[43] = 0000000000000000000000000000000000000000000000001110101101010010
# KERNEL: data of a[42] = 0000000000000000000000000000000000000000000000110100101101001000
# KERNEL: data of a[41] = 0000000000000000000000000000000000000000000000101110010111100100
# KERNEL: data of a[40] = 0000000000000000000000000000000000000000000000100101101011111111
# KERNEL: data of a[39] = 0000000000000000000000000000000000000000000000101010010000000010
# KERNEL: data of a[38] = 0000000000000000000000000000000000000000000000001011101011101011
# KERNEL: data of a[37] = 0000000000000000000000000000000000000000000001000011111001001011
# KERNEL: data of a[36] = 0000000000000000000000000000000000000000000000101001011100001001
# KERNEL: data of a[35] = 0000000000000000000000000000000000000000000000111001100010011000
# KERNEL: data of a[34] = 0000000000000000000000000000000000000000000000001010000111010010
# KERNEL: data of a[33] = 0000000000000000000000000000000000000000000001000001101101000100
# KERNEL: data of a[32] = 0000000000000000000000000000000000000000000000100111010101011010
# KERNEL: data of a[31] = 0000000000000000000000000000000000000000000000100101001100110010
# KERNEL: data of a[30] = 0000000000000000000000000000000000000000000000101010011001100010
# KERNEL: data of a[29] = 0000000000000000000000000000000000000000000000010111001111001101
# KERNEL: data of a[28] = 0000000000000000000000000000000000000000000000111110001101000101
# KERNEL: data of a[27] = 0000000000000000000000000000000000000000000000011000100101000011
# KERNEL: data of a[26] = 0000000000000000000000000000000000000000000000100101001100110110
# KERNEL: data of a[25] = 0000000000000000000000000000000000000000000001010111100110111001
# KERNEL: data of a[24] = 0000000000000000000000000000000000000000000000101101011000111001
# KERNEL: data of a[23] = 0000000000000000000000000000000000000000000001011100011010001011
# KERNEL: data of a[22] = 0000000000000000000000000000000000000000000000001111111100100001
# KERNEL: data of a[21] = 0000000000000000000000000000000000000000000000110110001101001010
# KERNEL: data of a[20] = 0000000000000000000000000000000000000000000000011111011011111011
# KERNEL: data of a[19] = 0000000000000000000000000000000000000000000000100011111100111000
# KERNEL: data of a[18] = 0000000000000000000000000000000000000000000000010110010100000110
# KERNEL: data of a[17] = 0000000000000000000000000000000000000000000000011011001100110011
# KERNEL: data of a[16] = 0000000000000000000000000000000000000000000001011010000100110011
# KERNEL: data of a[15] = 0000000000000000000000000000000000000000000000110110101001111011
# KERNEL: data of a[14] = 0000000000000000000000000000000000000000000001000010000100110001
# KERNEL: data of a[13] = 0000000000000000000000000000000000000000000001100011000010111001
# KERNEL: data of a[12] = 0000000000000000000000000000000000000000000000010000111001010110
# KERNEL: data of a[11] = 0000000000000000000000000000000000000000000000010001000110101000
# KERNEL: data of a[10] = 0000000000000000000000000000000000000000000000000111011111111100
# KERNEL: data of a[9] = 0000000000000000000000000000000000000000000000010100110111010111
# KERNEL: data of a[8] = 0000000000000000000000000000000000000000000000000101111101101001
# KERNEL: data of a[7] = 0000000000000000000000000000000000000000000001011111110110010111
# KERNEL: data of a[6] = 0000000000000000000000000000000000000000000000000000011011000001
# KERNEL: data of a[5] = 0000000000000000000000000000000000000000000000110011000110101000
# KERNEL: data of a[4] = 0000000000000000000000000000000000000000000001000110110011101010
# KERNEL: data of a[3] = 0000000000000000000000000000000000000000000000000010110001011110
# KERNEL: data of a[2] = 0000000000000000000000000000000000000000000001000101001001010100
# KERNEL: data of a[1] = 0000000000000000000000000000000000000000000000111111101110110110
# KERNEL: data of a[0] = 0000000000000000000000000000000000000000000000000011011101011111
# KERNEL: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.
