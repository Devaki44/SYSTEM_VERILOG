module code;
	int a;

	initial begin
		a= 32'b0101 ;
		$display(" %b",a);
	end
endmodule
