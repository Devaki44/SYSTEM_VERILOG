module repeat_loop;
  
  initial begin
    repeat(5)begin
      $display("BELIEVE YOURSELF");
    end
  end
endmodule



# KERNEL: BELIEVE YOURSELF
# KERNEL: BELIEVE YOURSELF
# KERNEL: BELIEVE YOURSELF
# KERNEL: BELIEVE YOURSELF
# KERNEL: BELIEVE YOURSELF
# KERNEL: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.
