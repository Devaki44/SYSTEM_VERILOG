//SAME FOR REG,LOGIC,BIT

module multi_dim_array;
  logic [3:0][1:0]a[7:0][3:0];
  
  initial begin
    
    foreach(a[i,j,k,l])begin
      
      a[i][j][k][l] = $urandom_range(0,256);
      
      $display("data of a[%0d][%0d][%0d][%0d] = %b",i,j,k,l,a[i][j][k][l]);
    end
  end
endmodule



# KERNEL: data of a[7][3][3][1] = 0
# KERNEL: data of a[7][3][3][0] = 1
# KERNEL: data of a[7][3][2][1] = 0
# KERNEL: data of a[7][3][2][0] = 0
# KERNEL: data of a[7][3][1][1] = 0
# KERNEL: data of a[7][3][1][0] = 0
# KERNEL: data of a[7][3][0][1] = 1
# KERNEL: data of a[7][3][0][0] = 0
# KERNEL: data of a[7][2][3][1] = 0
# KERNEL: data of a[7][2][3][0] = 1
# KERNEL: data of a[7][2][2][1] = 1
# KERNEL: data of a[7][2][2][0] = 1
# KERNEL: data of a[7][2][1][1] = 1
# KERNEL: data of a[7][2][1][0] = 1
# KERNEL: data of a[7][2][0][1] = 1
# KERNEL: data of a[7][2][0][0] = 1
# KERNEL: data of a[7][1][3][1] = 0
# KERNEL: data of a[7][1][3][0] = 1
# KERNEL: data of a[7][1][2][1] = 0
# KERNEL: data of a[7][1][2][0] = 0
# KERNEL: data of a[7][1][1][1] = 0
# KERNEL: data of a[7][1][1][0] = 0
# KERNEL: data of a[7][1][0][1] = 0
# KERNEL: data of a[7][1][0][0] = 1
# KERNEL: data of a[7][0][3][1] = 0
# KERNEL: data of a[7][0][3][0] = 0
# KERNEL: data of a[7][0][2][1] = 1
# KERNEL: data of a[7][0][2][0] = 0
# KERNEL: data of a[7][0][1][1] = 1
# KERNEL: data of a[7][0][1][0] = 0
# KERNEL: data of a[7][0][0][1] = 0
# KERNEL: data of a[7][0][0][0] = 0
# KERNEL: data of a[6][3][3][1] = 0
# KERNEL: data of a[6][3][3][0] = 0
# KERNEL: data of a[6][3][2][1] = 1
# KERNEL: data of a[6][3][2][0] = 1
# KERNEL: data of a[6][3][1][1] = 1
# KERNEL: data of a[6][3][1][0] = 0
# KERNEL: data of a[6][3][0][1] = 1
# KERNEL: data of a[6][3][0][0] = 0
# KERNEL: data of a[6][2][3][1] = 0
# KERNEL: data of a[6][2][3][0] = 1
# KERNEL: data of a[6][2][2][1] = 1
# KERNEL: data of a[6][2][2][0] = 0
# KERNEL: data of a[6][2][1][1] = 0
# KERNEL: data of a[6][2][1][0] = 1
# KERNEL: data of a[6][2][0][1] = 1
# KERNEL: data of a[6][2][0][0] = 1
# KERNEL: data of a[6][1][3][1] = 1
# KERNEL: data of a[6][1][3][0] = 1
# KERNEL: data of a[6][1][2][1] = 0
# KERNEL: data of a[6][1][2][0] = 0
# KERNEL: data of a[6][1][1][1] = 0
# KERNEL: data of a[6][1][1][0] = 1
# KERNEL: data of a[6][1][0][1] = 1
# KERNEL: data of a[6][1][0][0] = 1
# KERNEL: data of a[6][0][3][1] = 0
# KERNEL: data of a[6][0][3][0] = 1
# KERNEL: data of a[6][0][2][1] = 0
# KERNEL: data of a[6][0][2][0] = 0
# KERNEL: data of a[6][0][1][1] = 0
# KERNEL: data of a[6][0][1][0] = 1
# KERNEL: data of a[6][0][0][1] = 0
# KERNEL: data of a[6][0][0][0] = 1
# KERNEL: data of a[5][3][3][1] = 0
# KERNEL: data of a[5][3][3][0] = 1
# KERNEL: data of a[5][3][2][1] = 1
# KERNEL: data of a[5][3][2][0] = 0
# KERNEL: data of a[5][3][1][1] = 1
# KERNEL: data of a[5][3][1][0] = 0
# KERNEL: data of a[5][3][0][1] = 1
# KERNEL: data of a[5][3][0][0] = 0
# KERNEL: data of a[5][2][3][1] = 1
# KERNEL: data of a[5][2][3][0] = 1
# KERNEL: data of a[5][2][2][1] = 0
# KERNEL: data of a[5][2][2][0] = 1
# KERNEL: data of a[5][2][1][1] = 0
# KERNEL: data of a[5][2][1][0] = 0
# KERNEL: data of a[5][2][0][1] = 1
# KERNEL: data of a[5][2][0][0] = 0
# KERNEL: data of a[5][1][3][1] = 0
# KERNEL: data of a[5][1][3][0] = 0
# KERNEL: data of a[5][1][2][1] = 0
# KERNEL: data of a[5][1][2][0] = 1
# KERNEL: data of a[5][1][1][1] = 1
# KERNEL: data of a[5][1][1][0] = 0
# KERNEL: data of a[5][1][0][1] = 1
# KERNEL: data of a[5][1][0][0] = 0
# KERNEL: data of a[5][0][3][1] = 1
# KERNEL: data of a[5][0][3][0] = 0
# KERNEL: data of a[5][0][2][1] = 0
# KERNEL: data of a[5][0][2][0] = 0
# KERNEL: data of a[5][0][1][1] = 1
# KERNEL: data of a[5][0][1][0] = 0
# KERNEL: data of a[5][0][0][1] = 0
# KERNEL: data of a[5][0][0][0] = 1
# KERNEL: data of a[4][3][3][1] = 0
# KERNEL: data of a[4][3][3][0] = 1
# KERNEL: data of a[4][3][2][1] = 1
# KERNEL: data of a[4][3][2][0] = 0
# KERNEL: data of a[4][3][1][1] = 1
# KERNEL: data of a[4][3][1][0] = 0
# KERNEL: data of a[4][3][0][1] = 0
# KERNEL: data of a[4][3][0][0] = 0
# KERNEL: data of a[4][2][3][1] = 1
# KERNEL: data of a[4][2][3][0] = 0
# KERNEL: data of a[4][2][2][1] = 0
# KERNEL: data of a[4][2][2][0] = 1
# KERNEL: data of a[4][2][1][1] = 1
# KERNEL: data of a[4][2][1][0] = 0
# KERNEL: data of a[4][2][0][1] = 1
# KERNEL: data of a[4][2][0][0] = 1
# KERNEL: data of a[4][1][3][1] = 1
# KERNEL: data of a[4][1][3][0] = 1
# KERNEL: data of a[4][1][2][1] = 0
# KERNEL: data of a[4][1][2][0] = 0
# KERNEL: data of a[4][1][1][1] = 1
# KERNEL: data of a[4][1][1][0] = 1
# KERNEL: data of a[4][1][0][1] = 1
# KERNEL: data of a[4][1][0][0] = 0
# KERNEL: data of a[4][0][3][1] = 1
# KERNEL: data of a[4][0][3][0] = 0
# KERNEL: data of a[4][0][2][1] = 1
# KERNEL: data of a[4][0][2][0] = 0
# KERNEL: data of a[4][0][1][1] = 0
# KERNEL: data of a[4][0][1][0] = 0
# KERNEL: data of a[4][0][0][1] = 0
# KERNEL: data of a[4][0][0][0] = 0
# KERNEL: data of a[3][3][3][1] = 1
# KERNEL: data of a[3][3][3][0] = 1
# KERNEL: data of a[3][3][2][1] = 0
# KERNEL: data of a[3][3][2][0] = 0
# KERNEL: data of a[3][3][1][1] = 0
# KERNEL: data of a[3][3][1][0] = 1
# KERNEL: data of a[3][3][0][1] = 1
# KERNEL: data of a[3][3][0][0] = 0
# KERNEL: data of a[3][2][3][1] = 0
# KERNEL: data of a[3][2][3][0] = 0
# KERNEL: data of a[3][2][2][1] = 0
# KERNEL: data of a[3][2][2][0] = 0
# KERNEL: data of a[3][2][1][1] = 1
# KERNEL: data of a[3][2][1][0] = 1
# KERNEL: data of a[3][2][0][1] = 0
# KERNEL: data of a[3][2][0][0] = 0
# KERNEL: data of a[3][1][3][1] = 0
# KERNEL: data of a[3][1][3][0] = 1
# KERNEL: data of a[3][1][2][1] = 0
# KERNEL: data of a[3][1][2][0] = 0
# KERNEL: data of a[3][1][1][1] = 0
# KERNEL: data of a[3][1][1][0] = 1
# KERNEL: data of a[3][1][0][1] = 0
# KERNEL: data of a[3][1][0][0] = 1
# KERNEL: data of a[3][0][3][1] = 0
# KERNEL: data of a[3][0][3][0] = 1
# KERNEL: data of a[3][0][2][1] = 1
# KERNEL: data of a[3][0][2][0] = 1
# KERNEL: data of a[3][0][1][1] = 0
# KERNEL: data of a[3][0][1][0] = 0
# KERNEL: data of a[3][0][0][1] = 1
# KERNEL: data of a[3][0][0][0] = 0
# KERNEL: data of a[2][3][3][1] = 0
# KERNEL: data of a[2][3][3][0] = 0
# KERNEL: data of a[2][3][2][1] = 0
# KERNEL: data of a[2][3][2][0] = 0
# KERNEL: data of a[2][3][1][1] = 0
# KERNEL: data of a[2][3][1][0] = 0
# KERNEL: data of a[2][3][0][1] = 1
# KERNEL: data of a[2][3][0][0] = 0
# KERNEL: data of a[2][2][3][1] = 0
# KERNEL: data of a[2][2][3][0] = 0
# KERNEL: data of a[2][2][2][1] = 0
# KERNEL: data of a[2][2][2][0] = 1
# KERNEL: data of a[2][2][1][1] = 1
# KERNEL: data of a[2][2][1][0] = 1
# KERNEL: data of a[2][2][0][1] = 0
# KERNEL: data of a[2][2][0][0] = 0
# KERNEL: data of a[2][1][3][1] = 1
# KERNEL: data of a[2][1][3][0] = 0
# KERNEL: data of a[2][1][2][1] = 1
# KERNEL: data of a[2][1][2][0] = 0
# KERNEL: data of a[2][1][1][1] = 1
# KERNEL: data of a[2][1][1][0] = 1
# KERNEL: data of a[2][1][0][1] = 1
# KERNEL: data of a[2][1][0][0] = 1
# KERNEL: data of a[2][0][3][1] = 1
# KERNEL: data of a[2][0][3][0] = 1
# KERNEL: data of a[2][0][2][1] = 0
# KERNEL: data of a[2][0][2][0] = 1
# KERNEL: data of a[2][0][1][1] = 0
# KERNEL: data of a[2][0][1][0] = 1
# KERNEL: data of a[2][0][0][1] = 1
# KERNEL: data of a[2][0][0][0] = 0
# KERNEL: data of a[1][3][3][1] = 1
# KERNEL: data of a[1][3][3][0] = 1
# KERNEL: data of a[1][3][2][1] = 1
# KERNEL: data of a[1][3][2][0] = 1
# KERNEL: data of a[1][3][1][1] = 1
# KERNEL: data of a[1][3][1][0] = 1
# KERNEL: data of a[1][3][0][1] = 1
# KERNEL: data of a[1][3][0][0] = 0
# KERNEL: data of a[1][2][3][1] = 0
# KERNEL: data of a[1][2][3][0] = 1
# KERNEL: data of a[1][2][2][1] = 1
# KERNEL: data of a[1][2][2][0] = 0
# KERNEL: data of a[1][2][1][1] = 1
# KERNEL: data of a[1][2][1][0] = 0
# KERNEL: data of a[1][2][0][1] = 0
# KERNEL: data of a[1][2][0][0] = 0
# KERNEL: data of a[1][1][3][1] = 0
# KERNEL: data of a[1][1][3][0] = 0
# KERNEL: data of a[1][1][2][1] = 1
# KERNEL: data of a[1][1][2][0] = 0
# KERNEL: data of a[1][1][1][1] = 0
# KERNEL: data of a[1][1][1][0] = 1
# KERNEL: data of a[1][1][0][1] = 0
# KERNEL: data of a[1][1][0][0] = 1
# KERNEL: data of a[1][0][3][1] = 1
# KERNEL: data of a[1][0][3][0] = 0
# KERNEL: data of a[1][0][2][1] = 1
# KERNEL: data of a[1][0][2][0] = 1
# KERNEL: data of a[1][0][1][1] = 0
# KERNEL: data of a[1][0][1][0] = 1
# KERNEL: data of a[1][0][0][1] = 0
# KERNEL: data of a[1][0][0][0] = 0
# KERNEL: data of a[0][3][3][1] = 0
# KERNEL: data of a[0][3][3][0] = 1
# KERNEL: data of a[0][3][2][1] = 1
# KERNEL: data of a[0][3][2][0] = 1
# KERNEL: data of a[0][3][1][1] = 0
# KERNEL: data of a[0][3][1][0] = 0
# KERNEL: data of a[0][3][0][1] = 0
# KERNEL: data of a[0][3][0][0] = 1
# KERNEL: data of a[0][2][3][1] = 0
# KERNEL: data of a[0][2][3][0] = 1
# KERNEL: data of a[0][2][2][1] = 0
# KERNEL: data of a[0][2][2][0] = 1
# KERNEL: data of a[0][2][1][1] = 0
# KERNEL: data of a[0][2][1][0] = 0
# KERNEL: data of a[0][2][0][1] = 1
# KERNEL: data of a[0][2][0][0] = 0
# KERNEL: data of a[0][1][3][1] = 1
# KERNEL: data of a[0][1][3][0] = 0
# KERNEL: data of a[0][1][2][1] = 0
# KERNEL: data of a[0][1][2][0] = 0
# KERNEL: data of a[0][1][1][1] = 1
# KERNEL: data of a[0][1][1][0] = 0
# KERNEL: data of a[0][1][0][1] = 0
# KERNEL: data of a[0][1][0][0] = 0
# KERNEL: data of a[0][0][3][1] = 0
# KERNEL: data of a[0][0][3][0] = 1
# KERNEL: data of a[0][0][2][1] = 1
# KERNEL: data of a[0][0][2][0] = 1
# KERNEL: data of a[0][0][1][1] = 0
# KERNEL: data of a[0][0][1][0] = 0
# KERNEL: data of a[0][0][0][1] = 1
# KERNEL: data of a[0][0][0][0] = 1
# KERNEL: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.
